* Extracted by KLayout with SG13G2 LVS runset on : 10/04/2025 02:13

.SUBCKT Mixer5GHz GND ICC OSCN VCC OSCP IDC LOP IFP RFN LON VDC IFN RFP
M$1 GND ICC \$119878 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p
+ PS=133.9u PD=133.9u
M$21 GND ICC ICC GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p PS=133.9u
+ PD=133.9u
M$41 \$119878 OSCP OSCN GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$56 \$119878 OSCN OSCP GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$71 GND IDC \$590709 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p
+ PS=133.9u PD=133.9u
M$91 GND IDC IDC GND sg13_lv_nmos L=0.13u W=240u AS=47.4p AD=47.4p PS=267.8u
+ PD=267.8u
M$131 GND IDC \$590710 GND sg13_lv_nmos L=0.13u W=120u AS=23.7p AD=23.7p
+ PS=133.9u PD=133.9u
M$151 \$590709 LON LOP GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$166 \$590709 LOP LON GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p PS=102u
+ PD=102u
M$181 \$590710 IFP \$600001 GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p
+ PS=102u PD=102u
M$196 \$590710 IFN \$600002 GND sg13_lv_nmos L=0.13u W=90u AS=18p AD=18p
+ PS=102u PD=102u
M$211 \$600001 LOP RFP GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$221 \$600001 LON RFN GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$231 \$600002 LON RFP GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
M$241 \$600002 LOP RFN GND sg13_lv_nmos L=0.13u W=60u AS=12.3p AD=12.3p
+ PS=70.1u PD=70.1u
R$251 OSCP VCC rppd w=4.35u l=1.5u ps=0 b=0 m=1
R$252 OSCN VCC rppd w=4.35u l=1.5u ps=0 b=0 m=1
R$253 RFP VDC rppd w=4.5u l=3.2u ps=0 b=0 m=1
R$254 RFN VDC rppd w=4.5u l=3.2u ps=0 b=0 m=1
R$255 LON VDC rppd w=4.4u l=1.5u ps=0 b=0 m=1
R$256 LOP VDC rppd w=4.4u l=1.5u ps=0 b=0 m=1
C$257 VCC OSCP cap_cmim w=19.1u l=10.7u A=204.37p P=59.6u m=1
C$258 VCC OSCN cap_cmim w=19.1u l=10.7u A=204.37p P=59.6u m=1
C$259 VDC LOP cap_cmim w=11.745u l=9.445u A=110.931525p P=42.38u m=1
C$260 VDC LON cap_cmim w=11.745u l=9.445u A=110.931525p P=42.38u m=1
.ENDS Mixer5GHz
